grammar simple:extensions:list;

imports silver:langutil;
imports silver:langutil:pp;
imports simple:concretesyntax as cst;
imports simple:abstractsyntax;


terminal List 'List' lexer classes { KEYWORDS };

